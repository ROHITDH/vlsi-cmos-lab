*** SPICE deck for cell inverter{lay} from library VLSI_EXPERIMENTS
*** Created on Sat Mar 26, 2022 21:52:59
*** Last revised on Sat Mar 26, 2022 22:10:44
*** Written on Sat Mar 26, 2022 22:11:15 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: inverter{lay}
Mnmos@0 vout vin gnd gnd nmos L=0.4U W=2U AS=4.4P AD=2.4P PS=12.4U PD=6.4U
Mpmos@0 vout vin vdd vdd pmos L=0.4U W=2U AS=4.4P AD=2.4P PS=12.4U PD=6.4U

* Spice Code nodes in cell cell 'inverter{lay}'
vdd vdd 0 dc 5
vin vin 0 pulse 0 5 0 1n 1n 10n 20n
.tran 200n
.include C5_models.txt
.END
