*** SPICE deck for cell cs_amplifier{lay} from library VLSI_EXPERIMENTS
*** Created on Sun Mar 27, 2022 11:30:04
*** Last revised on Sun Mar 27, 2022 12:09:54
*** Written on Sun Mar 27, 2022 12:11:29 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: cs_amplifier{lay}
Mnmos@0 net@1 vbias gnd gnd nmos L=0.4U W=2U AS=5.6P AD=1.8P PS=14.4U PD=5.4U
Mnmos@1 gnd vin vout gnd nmos L=0.4U W=4U AS=3P AD=5.6P PS=7.4U PD=14.4U
Mpmos@0 vout net@1 vdd vdd pmos L=5U W=1U AS=1.7P AD=3P PS=5.4U PD=7.4U
Mpmos@2 vdd net@1 net@1 vdd pmos L=5U W=1U AS=1.8P AD=1.7P PS=5.4U PD=5.4U

* Spice Code nodes in cell cell 'cs_amplifier{lay}'
vdd vdd 0 dc 5
vbias vbias 0 dc 1.2
*dc analysis
*vin vin 0 dc 5
*.dc vin 0 5 0.1
*transient analysis
vin vin 0 ac sin(774.702m 5m 1k)
.tran 10m
*AC analysis
*vin vin 0 ac sin(offset 5m 1k)
*.ac DEC 100 100 10G
.include C5_models.txt
.END
