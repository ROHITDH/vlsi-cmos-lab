*** SPICE deck for cell cs_amplifier{sch} from library VLSI_EXPERIMENTS
*** Created on Sun Mar 27, 2022 09:38:53
*** Last revised on Sun Mar 27, 2022 09:59:41
*** Written on Sun Mar 27, 2022 10:10:46 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: cs_amplifier{sch}
Mnmos@0 net@6 vbias gnd gnd nmos L=0.4U W=2U
Mnmos@1 gnd vin vout gnd nmos L=0.4U W=4U
Mpmos@0 net@6 net@6 vdd vdd pmos L=5U W=1U
Mpmos@1 vdd net@6 vout vdd pmos L=5U W=1U

* Spice Code nodes in cell cell 'cs_amplifier{sch}'
vdd vdd 0 dc 5
vbias vbias 0 dc 1.2
*DC analysis
*----------------------------
*vin vin 0 dc 5
*.dc vin 0 5 0.1
*Transient Analysis
*-----------------------------
*V[name] n+ n- type sin(dc_offset amplitude frequency)
*vin vin 0 ac sin(0 1m 1k)
*.tran 100n
*AC analysis
*-----------------------------
vin vin 0 ac sin(774.615mV 1m 1k)
.ac DEC 100 100 10G
.include C5_models.txt
.END

